// Design Name:    basic_proc
// Module Name:    InstFetch 
// Project Name:   CSE141L
// Description:    instruction fetch (pgm ctr) for processor
//
// Revision:  2019.01.27
//
module ProgCtr #(parameter L=10) (
  input                Done, 
                       Reset,      // reset, init, etc. -- force PC to 0
                       Start,      // Signal to jump to next program; currently unused 
                       Clk,        // PC can change on pos. edges only
                       BranchRel,  // PC moves next line or line after 
							  Decision, // decides true or false for branches 
							  BranchAbs,  // jump to Target			
  input        [L-1:0] Target,     // jump ... "how high?"
  output logic [L-1:0] ProgCtr     // the program counter register itself
  );
  
   logic ever_start; 
   logic [3:0]first_start; 
   logic [3:0]second_start; 
   logic [3:0]third_start;

  // program counter can clear to 0, increment, or jump
  always_ff @(posedge Clk)	 begin           // or just always; always_ff is a linting construct
	if(Reset) begin
	    ProgCtr <= 0;				       // for first program; want different value for 2nd or 3rd
		ever_start <= '0;
		first_start <= '0;
		second_start <= '0;
		third_start <= '0;
	end else if(BranchAbs)	               // unconditional absolute jump
	  ProgCtr <= Target;			   //   how would you make it conditional and/or relative?
	else if(BranchRel) begin  // conditional relative jump
		if(Decision)
	  		ProgCtr <=  ProgCtr + 'b1;	   // if true go to the 2nd instruction 
		else 
			ProgCtr <= 	ProgCtr + 2'b10 ; 		// false so go to the next instruction 

    // else if (Ack) begin  

    //     // if (Start == 1) 
    //     //     ProgCtr <= ProgCtr+'b1;
    //     // else 
    //     ProgCtr <= ProgCtr;

    end else begin 

		if ( (first_start == '0) && (Start == '1) ) begin 
			first_start <= '1; 
		end else if ((first_start != '0) && (second_start == '0) && (Start == '1)) begin 
			second_start <= '1; 
		end else if ((first_start != '0) && (second_start != '0) && (third_start == '0) && (Start == '1)) begin 
			third_start <= '1;
		end

		if (Start == '1) begin 
			ever_start <= '1;
		end

		if (ever_start == '0) begin
			ProgCtr <= 0; 
		end else begin
			if (Start == '1) begin   
				ProgCtr <= ProgCtr; 
			end else if ( (first_start == '1) && (Start == '0) ) begin 
				ProgCtr <= 'b10; //prog 1 starts at 2
				first_start <= 'b10;
			end else if ( (second_start == '1) && (Start == '0) ) begin 
				ProgCtr <= 'b101000001; //prog 2 starts at 321
				second_start <= 'b10;
			end else if ( (third_start == '1) && (Start == '0) ) begin 
				ProgCtr <= 'b101000100;  //prog 3 starts at 324
				third_start <= 'b10;
			end else if (  (first_start == 'b10) || (second_start == 'b10) || (third_start == 'b10) ) 
                if (Done) 
                    ProgCtr <= ProgCtr; 
                else 
				    ProgCtr <= ProgCtr+'b1; //else just proceed like normal
		end

	end
  end //always end


endmodule


//added 2 dummy instructions in the start 
//added 2 dummy insns for prog2 
//changing jump for prog 3 to come back at the right instruction now










// 111101001
// 111101001
// 101010101
// 001101001
// 101001101
// 111000111
// 111000111
// 001000011
// 001000011
// 001000011
// 001000111
// 001000001
// 111011111
// 111011111
// 000011001
// 111001010
// 100001000
// 001000001
// 111001111
// 111001111
// 000001011
// 111001001
// 100001000
// 001000001
// 100011000
// 001000001
// 111011111
// 111011111
// 000011010
// 111010111
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010110 
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010101
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010100
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010011
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010010
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 111010001
// 100010000
// 001000001
// 111010111
// 111010111
// 000010011
// 100010000
// 111000111
// 111000111
// 111001111
// 111001111
// 001000011
// 001000011
// 001000011
// 001000111
// 001000001
// 000001000
// 101011000
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000010
// 001000001
// 100011000
// 000110011
// 111000111
// 111000111
// 000000001
// 101011000
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000010
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000111
// 001000001
// 100011000
// 111000111
// 111000111
// 000000001
// 101011000
// 001000001
// 101010000
// 011011010
// 001000111
// 001000001
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000111
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000111
// 101010000
// 011011010
// 001000111
// 001000001
// 100011000
// 111000111
// 111000111
// 000000001
// 101011000
// 001000111
// 101010000
// 011011010
// 001000111
// 101010000
// 011011010
// 001000111
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000111
// 101010000
// 011011010
// 001000001
// 101010000
// 011011010
// 001000010
// 100011000
// 111000111
// 111000111
// 000000001
// 001000010
// 001000111
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 001000001
// 101010000
// 011110010
// 011110011
// 001000111
// 100110000
// 111000111
// 111000111
// 010100000
// 001100001
// 000000001
// 101010000
// 010010100
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000001
// 101011000
// 010011100
// 000010011
// 111110001
// 001000010
// 001000001
// 101011000
// 010011100
// 000010011
// 111000111
// 111000111
// 000000001
// 001000010
// 001000111
// 001000001
// 101011000
// 010011100
// 111111001
// 001000001
// 101110000
// 010110100
// 000011110
// 111111001
// 001000001
// 101110000
// 010110100
// 000011110
// 111111001
// 001000111
// 001000001
// 101110000
// 010110100
// 000011110
// 111111001
// 111000111
// 111000111
// 010111000
// 000000001
// 001000110
// 001000111
// 101110000
// 010110100
// 000011110
// 111111001
// 001000111
// 001000001
// 101110000
// 010110100
// 000011110
// 111111001
// 001000001
// 101110000
// 010110100
// 000011110
// 111111001
// 001000001
// 101110000
// 010110100
// 000011110
// 001111101
// 001111110
// 001111010
// 001111001
// 111000111
// 111000111
// 000000111
// 001000111
// 000111101
// 100011111
// 001111001
// 100010111
// 111011111
// 111011111
// 000011101
// 001101001
// 110011100
// 110110000
// 111111111
// 111101001
// 111101011
// 111111111
// 111000111
// 111000111
// 010100000
// 010101000
// 010110000
// 010111000
// 010011000
// 001011011
// 001011011
// 001000000
// 101000000
// 111000011
// 111010111
// 111010111
// 010110010
// 000110100
// 101010011
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110001
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110010
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110011
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110100
// 111010011
// 111001111
// 111001111
// 000001011
// 001001001
// 101001001
// 111001111
// 000010001
// 110100010
// 001101001
// 101010011
// 111110101
// 111010011
// 111001111
// 111001111
// 000001011
// 001001001
// 101001001
// 111001110
// 000010001
// 110100010
// 001101001
// 101010011
// 111110110
// 111010011
// 111001111
// 111001111
// 000001011
// 001001001
// 101001001
// 111001101
// 000010001
// 110100010
// 001101001
// 101010011
// 111110111
// 111010011
// 111001111
// 111001111
// 000001011
// 001001001
// 101001001
// 111001100
// 000010001
// 110100010
// 001101001
// 001011001
// 111010111
// 111010111
// 000010110
// 111001111
// 111001111
// 000001100
// 110011001
// 001111001
// 110001101
// 110110011
// 111010111
// 111010111
// 010110010
// 000110100
// 101010011
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110001
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110010
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 101010011
// 111110011
// 111010011
// 110100010
// 001101001
// 110100010
// 001100001
// 111010111
// 111010111
// 000010110
// 111001111
// 111001111
// 000001100
// 110011001
// 001111001
// 001011100
// 001011001
// 100100011
// 001011001
// 100111011
// 001011001
// 100101011
// 111111111